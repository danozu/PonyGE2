library ieee;
        use ieee.std_logic_1164.all;
        
        entity tb is
        end tb;
        
        architecture test of tb is
        component ind1086708012
        port(d0: in std_ulogic; 
d1: in std_ulogic; 
d2: in std_ulogic; 
d3: in std_ulogic; 
d4: in std_ulogic; 
d5: in std_ulogic; 
d6: in std_ulogic; 
d7: in std_ulogic; 
a2: in std_ulogic; 
a1: in std_ulogic; 
a0: in std_ulogic; 
o: out std_ulogic); 
end component; 
signal d0, d1, d2, d3, d4, d5, d6, d7, a2, a1, a0, o: std_ulogic; 
begin 
ind1086708012ividual: ind1086708012  port map (d0 => d0, d1 => d1, d2 => d2, d3 => d3, d4 => d4, d5 => d5, d6 => d6, d7 => d7, a2 => a2, a1 => a1, a0 => a0, o => o); 
process begin 
d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '0';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '0';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '0';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '0';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '0';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '0';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '0';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '0';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '0';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '0';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '0';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

d0 <= '1';
d1 <= '1';
d2 <= '1';
d3 <= '1';
d4 <= '1';
d5 <= '1';
d6 <= '1';
d7 <= '1';
a2 <= '1';
a1 <= '1';
a0 <= '1';
wait for 1 ns; 
report std_ulogic'image(o) & CR;

	wait; 
	end process; 
end test;